************************************************************************
* Library Name: ICSN55H7RVT
* Cell Name:    OR2X1H7R
* View Name:    schematic
************************************************************************

.SUBCKT OR2X1H7R A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MMN2 net21 B VSS VSS nm1p2_svt_lp W=150n L=60n m=1
MMN0 net21 A VSS VSS nm1p2_svt_lp W=150n L=60n m=1
MMP2 net21 B net016 VDD pm1p2_svt_lp W=190n L=60n m=1
MMP1 net016 A VDD VDD pm1p2_svt_lp W=190n L=60n m=1
XXI4 net21 VDD VSS Y / INV pl=6e-08 pw=2.7e-07 nl=6e-08 nw=2.1e-07
.ENDS
